`timescale 1ns/1ps

module Booth_Multiplier_64_signed_tb();

    reg signed [63:0] a_i;
    reg signed [63:0] b_i;
    reg               clk;
    wire signed [127:0] result_o;

    Booth_Multiplier_64_signed uut (
        .a_i(a_i),
        .b_i(b_i),
        .clk(clk),
        .result_o(result_o)
    );

    always #5 clk = ~clk;
    initial begin
	    $dumpfile("Booth_Multiplier_64_signed_dump.vcd");
	    $dumpvars;
	    $dumpon;
        clk = 0;
	#10
        // Test case 1: 0 * 0
        a_i = 64'b0;
        b_i = 64'b0;
        #10;

        // Test case 2: 1 * 1
        a_i = 64'd1;
        b_i = 64'd1;
        #10;

        // Test case 3: -1 * -1
        a_i = -64'd1;
        b_i = -64'd1;
        #10;

        // Test case 4: 2^62 * 2^62
        a_i = 64'sd4611686018427387904;  // 2^62
        b_i = 64'sd4611686018427387904;  // 2^62
        #10;

        // Test case 5: -2^63 * 1
        a_i = -64'sd9223372036854775808;  // -2^63
        b_i = 64'd1;
        #10;

        // Test case 6: -2^63 * -1
        a_i = -64'sd9223372036854775808;  // -2^63
        b_i = -64'd1;
        #10;

        // Test case 7: -36 * 42
        a_i = -64'd36;
        b_i = 64'd42;
        #10;

        // Test case 8: 47 * 21
        a_i = 64'd47;
        b_i = 64'd21;
	#10

	//case 9: 55555*7777
	a_i = 64'd55555;
	b_i = 64'd77777;
	#10

	//case 10: 666666*333333
	a_i = 64'd666666;
	b_i = 64'd333333;
	#10
	
	//case 11: -987456321*205080080502
	a_i = -64'sd987456321;
	b_i = 64'd205080080502;
	#10

	//case 12: -9080706050*-40302010
	a_i = -64'sd9080706050;
	b_i = -64'sd40302010;
	#10
	
	//case 13: 987456321*-205080080502
	a_i = 64'd987456321;
	b_i = -64'sd205080080502;
	#10

	//case 14: 741852963*-55555555
	a_i = 64'd741852963;
	b_i = -64'sd55555555;
	#10

	//case 15: 74182963*-5555555
	a_i = 64'd74182963;
	b_i = -64'sd55555555;
	#10

	//case 16: 98987878*96967676
	a_i = 64'd98987878;
	b_i = 64'd96967676;
	#10

	//case 17: -7899851236547896*-2568
	a_i = -64'sd7899851236547896;
	b_i = -64'sd2568;
	#10

	//case 18: -147852365415245*158745698236547
	a_i = -64'sd147852365415245;
	b_i = 64'd158745698236547;
	#10

	//case 19: 789654123658745687*359874562587412568
	a_i = 64'd789654123658745687;
	b_i = 64'd359874562587412568;
	#10
	
	//case 20: -89654123658745687*-59874562587412568
	a_i = -64'sd89654123658745687;
	b_i = -64'sd59874562587412568;
	#10

        #30;
	$dumpoff;
	$dumpflush;
        $finish;  
    end

endmodule